* W:\TCO\pract_7\F_2.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 08 08:59:59 2018



** Analysis setup **
.tran 0ns 1u
.LIB "W:\TCO\pract_7\NAND_1.lib"
.STMLIB "F_2.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "F_2.net"
.INC "F_2.als"


.probe


.END
