* W:\TCO\pract_4\ejer_1.sch

* Schematics Version 9.1 - Web Update 1
* Tue Mar 06 09:03:02 2018



** Analysis setup **
.DC LIN V_VGS 0 5 0.1 
.OP 
.LIB "W:\TCO\pract_4\ejer_1.lib"
.STMLIB "ejer_1.stl"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "ejer_1.net"
.INC "ejer_1.als"


.probe


.END
