* W:\TCO\pract_7\NAND_1.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 08 08:43:46 2018



** Analysis setup **
.OP 
.LIB "W:\TCO\pract_7\NAND_1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NAND_1.net"
.INC "NAND_1.als"


.probe


.END
